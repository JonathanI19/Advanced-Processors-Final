module ALU_control(ALU_op, instruction, out);

    // I/O
    input [1:0] ALU_op;
    input 





endmodule:  ALU_control